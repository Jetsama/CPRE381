
library IEEE;
use IEEE.std_logic_1164.all;

entity tb_regFile is
  generic(gCLK_HPER   : time := 50 ns);
end tb_regFile;

architecture behavior of tb_regFile is
  
  -- Calculate the clock period as twice the half-period
  constant cCLK_PER  : time := gCLK_HPER * 2;


	component regFile is
  	generic(N : integer := 32); -- Generic of type integer for input/output data width. Default value is 32.
  	port(i_SR0          : in std_logic_vector(5-1 downto 0);
	i_SR1          : in std_logic_vector(5-1 downto 0);
       i_SW         : in std_logic_vector(5-1 downto 0);
	i_D          : in std_logic_vector(N-1 downto 0);

	i_CLK         : in std_logic;
	i_RST         : in std_logic;

       o_R0          : out std_logic_vector(N-1 downto 0);
	o_R1          : out std_logic_vector(N-1 downto 0));
	  end component;


  -- Temporary signals to connect to the dff component.
  signal s_CLK, s_RST, s_WE  : std_logic;
signal s_SR0, s_SR1,s_SW : std_logic_vector(5-1 downto 0);
  signal s_R0, s_R1,s_D : std_logic_vector(32-1 downto 0);

begin

  DUT: regFile 
  port map(i_CLK => s_CLK, 
           i_RST => s_RST,
           i_SW  => s_SW,
           i_SR1   => s_SR1,
		i_SR0   => s_SR0,
		i_D   => s_D,
		o_R0   => s_R0,
           o_R1   => s_R1);

  -- This process sets the clock value (low for gCLK_HPER, then high
  -- for gCLK_HPER). Absent a "wait" command, processes restart 
  -- at the beginning once they have reached the final statement.
  P_CLK: process
  begin
    s_CLK <= '0';
    wait for gCLK_HPER;
    s_CLK <= '1';
    wait for gCLK_HPER;
  end process;
  
  -- Testbench process  
  P_TB: process
  begin

s_SW  <= "00000";
	s_SR0 <= "00000";
	s_SR1  <= "00000";
s_D <= x"00000100";
    wait for cCLK_PER;

    -- Store '1'
    s_RST <= '0';
    s_WE  <= '1';
    s_D   <= x"00000001";
    wait for cCLK_PER;  

    -- Keep '1'

    s_D   <= x"00000000";
    wait for cCLK_PER;  

    -- Store '5'    
	s_SR0 <= "00001";
	s_SW  <= "00001";
	s_SR1  <= "00000";
    s_D   <= x"00000101";
    wait for cCLK_PER;  

    -- Keep '0'
	s_SR0 <= "00001";
	s_SW  <= "00011";
	s_SR1  <= "00000";
    s_D   <= x"00000111";
    s_D   <= x"00000001";
    wait for cCLK_PER;  
s_SR0 <= "00001";
	s_SW  <= "00011";	s_SR1  <= "00000";
    s_D   <= x"00000111";
    s_D   <= x"00000001";
    wait for cCLK_PER;  
    wait;
  end process;
  
end behavior;